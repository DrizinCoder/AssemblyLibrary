module Buffer(

	input [16:0] Numbers,
	output [7:0] element

);


endmodule
