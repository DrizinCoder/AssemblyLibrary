module AXI_Slave_Interface();


endmodule
