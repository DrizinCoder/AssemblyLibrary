module Sum(
	
	input [7:0] Num1,
	input [7:0] Num2,
	output [7:0] res
	
);

	assign res = Num1 + Num2;

endmodule
